module step_sequencer(
    // Inputs
    input wire	      CLOCK_50,
    input wire	[3:0] KEY,

    // Outputs
    output wire [6:0] HEX0,
    output wire [6:0] HEX1,
    output wire [6:0] HEX2,
    output wire [6:0] HEX3,
    output wire [6:0] HEX4,
    output wire [6:0] HEX5,
    output wire [9:0] LEDR,
	 
	output wire  	  AUD_XCK,
	output wire 	  AUD_DACDAT,

	output wire   	  FPGA_I2C_SCLK,
	output wire 	  DAC_I2C_SCLK, // PIN_Y17,  GPIO_0[1]
	output wire 	  DAC_I2C_A0,   // PIN_AD17, GPIO_0[2]

	output wire [7:0] VGA_R,
    output wire [7:0] VGA_G,
    output wire [7:0] VGA_B,
    output wire       VGA_HS,
    output wire       VGA_VS,
    output wire       VGA_BLANK_N,
    output wire       VGA_SYNC_N,
    output wire       VGA_CLK,  
	 
	// Bidirectionals
	inout wire   	  AUD_BCLK,
	inout wire 	      AUD_ADCLRCK,
	inout wire 	      AUD_DACLRCK,

	inout wire   	  FPGA_I2C_SDAT,
	inout wire 	      DAC_I2C_SDAT, // PIN_AC18, GPIO_0[0]
	 
	inout wire 	      PS2_CLK,
    inout wire 		  PS2_DAT
);
	 
	// Internal wires
	wire        nReset;
	wire [11:0] select_val;
	 
	wire        start_playback;
	wire [6:0]  loops_val;
	wire [9:0]  bpm_val;
	wire [3:0]  dir_val;
	wire 		cmd_val;
	wire        bpm_step;  // pulse generated by bpm
	wire   	    play_en;   // play while this signal is high
	 
	 
	// Combinational logic
	assign nReset = KEY[0];

	// Start pulse
	reg start_prev;
   	always@(posedge CLOCK_50, negedge nReset)
   	begin   
    	if (!nReset)
    	begin
        	start_prev <= 0;
    	end
    	else
    	begin
        	start_prev <= start_playback;
    	end
   	end

   wire start_pulse = (start_playback && start_prev != 1);
	
	audio_interface A1 (
		// Inputs
		.CLOCK_50      (CLOCK_50),
		.nStart        (~start_pulse), // Start playback
		.nReset        (nReset),          // Reset
		.Select        (select_val),	  // Tone select
		.Loops         (loops_val),       // Number of playback loops
		.BPM           (bpm_val),         // Beats per minute
		
		// Bidirectionals
		.AUD_BCLK      (AUD_BCLK),
		.AUD_ADCLRCK   (AUD_ADCLRCK ),
		.AUD_DACLRCK   (AUD_DACLRCK ),

		.FPGA_I2C_SDAT (FPGA_I2C_SDAT),
		.DAC_I2C_SDAT  (DAC_I2C_SDAT),    // PIN_AC18, GPIO_0[0]

		// Outputs
		.bpm_step 	   (bpm_step),
		.play_en	   (play_en),

		.AUD_XCK       (AUD_XCK),
		.AUD_DACDAT    (AUD_DACDAT),

		.FPGA_I2C_SCLK (FPGA_I2C_SCLK),
		.DAC_I2C_SCLK  (DAC_I2C_SCLK ),   // PIN_Y17,  GPIO_0[1]
		.DAC_I2C_A0    (DAC_I2C_A0)       // PIN_AD17, GPIO_0[2]
	);
	
	input_interface I1 (
		// Inputs
		.CLOCK_50  (CLOCK_50),
		.nReset    (nReset),
		.play_en   (play_en),

		// Outputs
		.HEX0 	   (HEX0),
		.HEX1 	   (HEX1),
		.HEX2 	   (HEX2),
		.HEX3 	   (HEX3),
		.HEX4 	   (HEX4),
		.HEX5 	   (HEX5),
		.LEDR 	   (LEDR),

		.BPM	   (bpm_val),
		.Loops     (loops_val),
		.Direction (dir_val),
		.Command   (cmd_val),
		.Start     (start_playback),

		// Bidirectionals
		.PS2_CLK   (PS2_CLK),
		.PS2_DAT   (PS2_DAT)
	);

	display_interface D1 (
		.CLOCK_50    (CLOCK_50),
		.nReset      (nReset),

		.Direction   (dir_val),
		.Command     (cmd_val),
		.play_en     (play_en),   // Playback enable
        .bpm_step    (bpm_step),  // BPM pulse
		.select_note (select_val),

		.VGA_R       (VGA_R),
        .VGA_G       (VGA_G),
        .VGA_B       (VGA_B),
        .VGA_HS      (VGA_HS),
        .VGA_VS      (VGA_VS),
        .VGA_BLANK_N (VGA_BLANK_N),
        .VGA_SYNC_N  (VGA_SYNC_N),
        .VGA_CLK     (VGA_CLK)	
	);

endmodule


