module BPM_counter (Clock, nStart, BPM, Step);
	input Clock, nStart;
   input [31:0] BPM; // Max 511 BPM [8:0]
	output reg Step;

   reg [31:0] Q;
   reg [63:0] target; 
   always@(posedge Clock, negedge nStart)
   begin
		// target = freq_clock * 60/BPM
      target = (64'd50_000_000 * 60) / BPM;
      if (!nStart)
      begin
          Step <= 0;
          Q <= 0;
      end
      else if (!BPM)
      begin
          Step <= 0;
          Q <= 0;
      end
      else if (Q == target)
      begin
          Q <= 0;
          Step <= 1;
      end       
      else
      begin
          Q <= Q + 1;
          Step <= 0;
      end 
    end
endmodule