module loop_counter (nReset, nStart, Step, Loops, Play);
    input nReset, nStart, Step;
    input [6:0] Loops; // Max 255 Loops
    output reg Play;

    reg [11:0] Q;
    reg [11:0] total_steps;
    reg done;
	 reg [6:0] Loops_latched;
	 
	 always@(posedge Step, negedge nReset, negedge nStart)
	 begin
	   if (!nReset)
		begin
			done          <= 1;
			Play 			  <= 0;
			Q             <= 0;
	   end
		else if (!nStart)
		begin
			Loops_latched <= Loops;
			done          <= 0;
			Play 			  <= 1;
			Q             <= 0;
			total_steps   <= Loops * 16;
	   end
		else if (Loops_latched == 0 && !done)
			Play <= 1;
		else if (!done)
		begin
			if (Q == total_steps - 1)
			begin
				done   <= 1;
				Play   <= 0;
			end
			else
			begin
				Play <= 1;
				Q    <= Q + 1;
			end
		end
		else
		begin
			done   <= 1;
			Play   <= 0;
		end
	 end
	 
endmodule