`default_nettype none
module vga_display (
    input  wire        CLOCK_50,
    input  wire        nReset,
    input  wire        state,        // 1 = white, 0 = blue
    input  wire        draw_enable,  // 1-cycle start pulse

    input  wire [9:0]  X,            // center or reference point
    input  wire [8:0]  Y,

    output reg         drawing,      // 1 while drawing 30x30 block

    output wire [9:0]  VGA_X,
    output wire [8:0]  VGA_Y, 
    output wire [23:0] VGA_COLOR, 
    output wire        plot
);

    // Internal registers
    reg [9:0] current_x;
    reg [8:0] current_y;
    reg       write;

    reg [1:0] current_state, next_state;

    reg [4:0] dx; 
    reg [4:0] dy;  

    reg [8:0] color;  
    wire      VGA_SYNC;

    // State parameters
    localparam IDLE = 2'b01,
               DRAW = 2'b10;

    always @(posedge CLOCK_50 or negedge nReset) begin
        if (!nReset) 
        begin
            color <= 9'd0;
        end 
        else if (draw_enable) 
        begin
            color <= state ? 9'h1FF : 9'd7;
        end
    end

    // State logic
    always @(*) begin
        if (!VGA_SYNC)
            next_state = IDLE;
        else begin
            case (current_state)
                IDLE:
                    next_state = draw_enable ? DRAW : IDLE;
                DRAW:
                    next_state = (!drawing) ? IDLE : DRAW;

                default:
                    next_state = IDLE;
            endcase
        end
    end
    
    // Drawing logic
    always @(posedge CLOCK_50 or negedge nReset) begin
        if (!nReset) 
        begin
            current_state <= IDLE;
            drawing       <= 0;
            write         <= 0;
            current_x     <= 0;
            current_y     <= 0;
            dx            <= 0;
            dy            <= 0;
        end 
        else if (!VGA_SYNC) 
        begin
            current_state <= IDLE;
            drawing       <= 0;
            write         <= 0;
            dx            <= 0;
            dy            <= 0;
        end 
        else 
        begin
            current_state <= next_state;
            case (next_state)
                IDLE: 
                begin
                    drawing   <= 0;
                    write     <= 0;
                    dx        <= 0;
                    dy        <= 0;
                   
                    current_x <= X;
                    current_y <= Y;
                end
                DRAW: 
                begin
                    drawing <= 1;
                    write   <= 1;

                    current_x <= X + dx;
                    current_y <= Y + dy;

                    if (dx < 30) begin
                        dx <= dx + 1;
                    end else begin
                        dx <= 0;
                        if (dy < 30)
                            dy <= dy + 1;
                        else
                            drawing <= 0; 
                    end
                end
            endcase
        end
    end

    // VGA adapter
    `define VGA_MEMORY
    vga_adapter VGA (
        .resetn    (nReset),
        .clock     (CLOCK_50),
        .color     (color),
        .x         (current_x),
        .y         (current_y),
        .write     (write),

        .VGA_X     (VGA_X),
        .VGA_Y     (VGA_Y),
        .VGA_COLOR (VGA_COLOR),
        .VGA_SYNC  (VGA_SYNC),
        .plot      (plot)
    );
    defparam VGA.RESOLUTION       = "640x480";
    defparam VGA.BACKGROUND_IMAGE = "./MIF/grid.mif";
    defparam VGA.COLOR_DEPTH      = 9;

endmodule