module step_sequencer (
    // Inputs
    input wire	      CLOCK_50,
    input wire	[2:0] KEY,

    // Outputs
    output wire [6:0] HEX0,
    output wire [6:0] HEX1,
    output wire [6:0] HEX2,
    output wire [6:0] HEX3,
    output wire [6:0] HEX4,
    output wire [6:0] HEX5,
    output wire [9:0] LEDR,
	 
	input wire  [8:0] sim_data,
	input wire        sim_data_en
);
	// Sim wires
	wire [9:0]  VGA_X;
    wire [8:0]  VGA_Y;
    wire [23:0] VGA_COLOR;
    wire        plot;   

	wire        AUD_XCK;
	wire 	    AUD_DACDAT;

	wire   	    FPGA_I2C_SCLK;
	wire 	    DAC_I2C_SCLK; // PIN_Y17,  GPIO_0[1]
	wire 	    DAC_I2C_A0;  // PIN_AD17, GPIO_0[2]
	 
	// Bidirectionals
	wire   	    AUD_BCLK;
	wire 	    AUD_ADCLRCK;
	wire 	    AUD_DACLRCK;

	wire   	    FPGA_I2C_SDAT;
	wire 	    DAC_I2C_SDAT; // PIN_AC18, GPIO_0[0]
	 
	// Internal wires
	wire        nReset;
	wire [11:0] select_val;
	 
	wire        start_playback;
	wire [6:0]  loops_val;
	wire [9:0]  bpm_val;
	wire [3:0]  dir_val;
	wire 		cmd_val;
	wire        bpm_step;  // pulse generated by bpm
	wire   	    play_en;   // play while this signal is high
	 
	 
	// Combinational logic
	assign nReset = KEY[0];
	
	audio_interface A1 (
		// Inputs
		.CLOCK_50      (CLOCK_50),
		.nStart        (~start_playback), // Start playback
		.nReset        (nReset),          // Reset
		.Select        (select_val),	  // Tone select
		.Loops         (loops_val),       // Number of playback loops
		.BPM           (bpm_val),         // Beats per minute
		
		// Bidirectionals
		.AUD_BCLK      (AUD_BCLK),
		.AUD_ADCLRCK   (AUD_ADCLRCK ),
		.AUD_DACLRCK   (AUD_DACLRCK ),

		.FPGA_I2C_SDAT (FPGA_I2C_SDAT),
		.DAC_I2C_SDAT  (DAC_I2C_SDAT),    // PIN_AC18, GPIO_0[0]

		// Outputs
		.bpm_step 	   (bpm_step),
		.play_en	   (play_en),

		.AUD_XCK       (AUD_XCK),
		.AUD_DACDAT    (AUD_DACDAT),

		.FPGA_I2C_SCLK (FPGA_I2C_SCLK),
		.DAC_I2C_SCLK  (DAC_I2C_SCLK ),   // PIN_Y17,  GPIO_0[1]
		.DAC_I2C_A0    (DAC_I2C_A0)       // PIN_AD17, GPIO_0[2]
	);
	
	input_interface I1 (
		// Inputs
		.CLOCK_50  (CLOCK_50),
		.nReset    (nReset),
		.play_en   (play_en),

		// Outputs
		.HEX0 	   (HEX0),
		.HEX1 	   (HEX1),
		.HEX2 	   (HEX2),
		.HEX3 	   (HEX3),
		.HEX4 	   (HEX4),
		.HEX5 	   (HEX5),
		.LEDR 	   (LEDR),

		.BPM	   (bpm_val),
		.Loops     (loops_val),
		.Direction (dir_val),
		.Command   (cmd_val),
		.Start     (start_playback),

		// Bidirectionals
		.sim_data_en (sim_data_en),
		.sim_data    (sim_data)
	);

	display_interface D1 (
		.CLOCK_50 (CLOCK_50),
		.nReset   (nReset),

		.Direction (dir_val),
		.Command   (cmd_val),
		.play_en   (play_en),   // Playback enable
        .bpm_step  (bpm_step),  // BPM pulse
		.select_note (select_val),

        .VGA_X     (VGA_X),
        .VGA_Y     (VGA_Y),
        .VGA_COLOR (VGA_COLOR),
        .plot      (plot)
	);

endmodule


